library ieee_proposed;  use ieee_proposed.electrical_systems.all;
                        
entity inline_18a is

end entity inline_18a;


architecture test of inline_18a is

begin

  process is
  begin

    -- code from book

    break;

    -- end code from book

    wait;
  end process;

end architecture test;
