library ieee_proposed;
use ieee_proposed.electrical_systems.all;
use ieee_proposed.mechanical_systems.all;
                        
entity inline_01a is

end entity inline_01a;


architecture test of inline_01a is

  -- code from book

  alias ground is electrical_ref;

  --

  alias anchor is translational_ref;

  -- end code from book

begin
end architecture test;
