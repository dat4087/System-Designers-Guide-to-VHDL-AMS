entity inline_14a is

end entity inline_14a;


----------------------------------------------------------------


architecture test of inline_14a is

  -- code from book:

  type array3 is array (10 downto 1) of real tolerance "default";

  quantity a3 : array3;

  -- end of code from book
  
begin
end architecture test;
