package inline_08 is

  -- code from book

  procedure uniform ( variable seed1, seed2 : inout positive;
                      variable x : out real);

  -- end code from book

end package inline_08;
