entity top_level is
end entity top_level;
