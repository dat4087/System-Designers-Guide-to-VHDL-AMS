package pk_chap5 is

  subtype word is integer;

end package pk_chap5;
