entity inline_04d is

end entity inline_04d;


----------------------------------------------------------------


library ieee;

architecture test of inline_04d is
begin


  block_3_c : block is

    -- code from book:

    use ieee.std_logic_1164.all;

    -- end of code from book

  begin
  end block block_3_c;


end architecture test;
