entity ent is

end entity ent;

architecture sample of ent is

  constant pi : real := 3.14159;

begin

  process is
    variable counter : integer;
  begin
    -- . . .         --  statements using pi and counter
  end process;

end architecture sample;
