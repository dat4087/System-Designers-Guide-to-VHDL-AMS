entity inline_04a is

end entity inline_04a;


----------------------------------------------------------------


library ieee_proposed;

architecture test of inline_04a is
begin


  block_3_c : block is

    -- code from book:

    use ieee_proposed.electrical_systems.all;

    -- end of code from book

  begin
  end block block_3_c;


end architecture test;
