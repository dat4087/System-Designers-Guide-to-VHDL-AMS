package int_types is

  type small_int is range 0 to 255;

end package int_types;
