entity inline_02a is

end entity inline_02a;


----------------------------------------------------------------


library wasp_lib;

-- code from book:

use wasp_lib.all;

-- end of code from book


architecture test of inline_02a is
begin

end architecture test;
