entity controller is
end entity controller;


-- code from book

architecture instrumented of controller is

  shared variable operation_count : natural := 0;
  -- . . .

begin
  -- . . .
end architecture instrumented;

-- end code from book
