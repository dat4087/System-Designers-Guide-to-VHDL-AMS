use work.int_types.all;

entity small_adder is
  port ( a, b : in small_int;  s : out small_int );
end entity small_adder;
